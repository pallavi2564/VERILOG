module not(
  input a;
  output y;)
  assign y=~a;
endmodule
